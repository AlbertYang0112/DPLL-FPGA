`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    23:05:55 05/05/2018 
// Design Name:    
// Module Name:    DPLL 
// Project Name:   DPLL-FPGA
// Target Devices: XC6SLX9-2FTG256
// Tool versions: 
// Description:     The digital phase lock loop.
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module DPLL(
    input baseClockInput,
    input oscInput,
    output dpllOutput
    );


endmodule
